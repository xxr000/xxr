module top;
	initial begin
		$display("XXR");
	end
endmodule
